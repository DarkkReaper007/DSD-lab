`include "L44.v"

`timescale 1ns / 1ns

module L44_tb;

    reg [15:0] A;
    wire [3:0] Y;

    // Instantiate the 16-to-4 priority encoder
    L44 uut (
        A,
        Y
    );

    initial begin
        $dumpfile("L44_tb.vcd");
        $dumpvars(0, L44_tb);

        A = 16'b0000000000000000; #10;
        A = 16'b0000000000000001; #10;
        A = 16'b0000000000000010; #10;
        A = 16'b0000000000000100; #10;
        A = 16'b0000000000001000; #10;
        A = 16'b0000000000010000; #10;
        A = 16'b0000000000100000; #10;
        A = 16'b0000000001000000; #10;
        A = 16'b0000000010000000; #10;
        A = 16'b0000000100000000; #10;
        A = 16'b0000001000000000; #10;
        A = 16'b0000010000000000; #10;
        A = 16'b0000100000000000; #10;
        A = 16'b0001000000000000; #10;
        A = 16'b0010000000000000; #10;
        A = 16'b0100000000000000; #10;
        A = 16'b1000000000000000; #10;

        $display("Test Complete");
        $finish;
    end

endmodule

